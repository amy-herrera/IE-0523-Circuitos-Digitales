localparam [9:0] K28_0_rd_plus  = 10'b1100001011;
localparam [9:0] K28_0_rd_minus = 10'b0011110100;

localparam [9:0] K28_1_rd_plus  = 10'b1100000110;
localparam [9:0] K28_1_rd_minus = 10'b0011111001;

localparam [9:0] K28_2_rd_plus  = 10'b1100001010;
localparam [9:0] K28_2_rd_minus = 10'b0011110101;

localparam [9:0] K28_3_rd_plus  = 10'b1100001100;
localparam [9:0] K28_3_rd_minus = 10'b0011110011;

localparam [9:0] K28_4_rd_plus  = 10'b1100001101;
localparam [9:0] K28_4_rd_minus = 10'b0011110010;

localparam [9:0] K28_5_rd_plus  = 10'b1100000101;
localparam [9:0] K28_5_rd_minus = 10'b0011111010;

localparam [9:0] K28_6_rd_plus  = 10'b1100001001;
localparam [9:0] K28_6_rd_minus = 10'b0011110110;

localparam [9:0] K28_7_rd_plus  = 10'b1100000111;
localparam [9:0] K28_7_rd_minus = 10'b0011111000;

localparam [9:0] K23_7_rd_plus  = 10'b0001010111;
localparam [9:0] K23_7_rd_minus = 10'b1110101000;

localparam [9:0] K27_7_rd_plus  = 10'b0010010111;
localparam [9:0] K27_7_rd_minus = 10'b1101101000;

localparam [9:0] K29_7_rd_plus  = 10'b0100010111;
localparam [9:0] K29_7_rd_minus = 10'b1011101000;

localparam [9:0] K30_7_rd_plus  = 10'b1000010111;
localparam [9:0] K30_7_rd_minus = 10'b0111101000;

localparam [9:0] D0_0_rd_plus   = 10'b0110001011;
localparam [9:0] D0_0_rd_minus  = 10'b1001110100;

localparam [9:0] D1_0_rd_plus   = 10'b1000101011;
localparam [9:0] D1_0_rd_minus  = 10'b0111010100;

localparam [9:0] D2_0_rd_plus   = 10'b0100101011;
localparam [9:0] D2_0_rd_minus  = 10'b1011010100;

localparam [9:0] D3_0_rd_plus   = 10'b1100010100;
localparam [9:0] D3_0_rd_minus  = 10'b1100011011;

localparam [9:0] D4_0_rd_plus   = 10'b0010101011;
localparam [9:0] D4_0_rd_minus  = 10'b1101010100;

localparam [9:0] D5_0_rd_plus   = 10'b1010010100;
localparam [9:0] D5_0_rd_minus  = 10'b1010011011;

localparam [9:0] D6_0_rd_plus   = 10'b0110010100;
localparam [9:0] D6_0_rd_minus  = 10'b0110011011;

localparam [9:0] D7_0_rd_plus   = 10'b0001110100;
localparam [9:0] D7_0_rd_minus  = 10'b1110001011;

localparam [9:0] D8_0_rd_plus   = 10'b0001101011;
localparam [9:0] D8_0_rd_minus  = 10'b1110010100;

localparam [9:0] D5_6_rd_plus   = 10'b1010010110;
localparam [9:0] D5_6_rd_minus  = 10'b1010010110;

localparam [9:0] D16_2_rd_plus  = 10'b1001000101;
localparam [9:0] D16_2_rd_minus = 10'b0110110101;
